-- nios.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios is
	port (
		clk_clk                  : in  std_logic                     := '0'; --                 clk.clk
		gpio_export              : out std_logic_vector(31 downto 0);        --                gpio.export
		reset_reset_n            : in  std_logic                     := '0'; --               reset.reset_n
		spi_eeprom_external_MISO : in  std_logic                     := '0'; -- spi_eeprom_external.MISO
		spi_eeprom_external_MOSI : out std_logic;                            --                    .MOSI
		spi_eeprom_external_SCLK : out std_logic;                            --                    .SCLK
		spi_eeprom_external_SS_n : out std_logic;                            --                    .SS_n
		spi_enet_external_MISO   : in  std_logic                     := '0'; --   spi_enet_external.MISO
		spi_enet_external_MOSI   : out std_logic;                            --                    .MOSI
		spi_enet_external_SCLK   : out std_logic;                            --                    .SCLK
		spi_enet_external_SS_n   : out std_logic                             --                    .SS_n
	);
end entity nios;

architecture rtl of nios is
	component nios_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(15 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component nios_CPU;

	component nios_GPIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component nios_GPIO;

	component nios_RAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component nios_RAM;

	component nios_ROM is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			debugaccess : in  std_logic                     := 'X';             -- debugaccess
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component nios_ROM;

	component nios_SPI_EEPROM is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component nios_SPI_EEPROM;

	component nios_SPI_ENET is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component nios_SPI_ENET;

	component nios_SystemTick is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_SystemTick;

	component nios_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_jtag_uart_0;

	component nios_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest               : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                      : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_write                     : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess               : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address            : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest        : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read               : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_debug_mem_slave_address               : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write                 : out std_logic;                                        -- write
			CPU_debug_mem_slave_read                  : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess           : out std_logic;                                        -- debugaccess
			GPIO_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			GPIO_s1_write                             : out std_logic;                                        -- write
			GPIO_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			GPIO_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			GPIO_s1_chipselect                        : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			RAM_s1_address                            : out std_logic_vector(10 downto 0);                    -- address
			RAM_s1_write                              : out std_logic;                                        -- write
			RAM_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RAM_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			RAM_s1_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			RAM_s1_chipselect                         : out std_logic;                                        -- chipselect
			RAM_s1_clken                              : out std_logic;                                        -- clken
			ROM_s1_address                            : out std_logic_vector(12 downto 0);                    -- address
			ROM_s1_write                              : out std_logic;                                        -- write
			ROM_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ROM_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			ROM_s1_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			ROM_s1_chipselect                         : out std_logic;                                        -- chipselect
			ROM_s1_clken                              : out std_logic;                                        -- clken
			ROM_s1_debugaccess                        : out std_logic;                                        -- debugaccess
			SPI_EEPROM_spi_control_port_address       : out std_logic_vector(2 downto 0);                     -- address
			SPI_EEPROM_spi_control_port_write         : out std_logic;                                        -- write
			SPI_EEPROM_spi_control_port_read          : out std_logic;                                        -- read
			SPI_EEPROM_spi_control_port_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SPI_EEPROM_spi_control_port_writedata     : out std_logic_vector(15 downto 0);                    -- writedata
			SPI_EEPROM_spi_control_port_chipselect    : out std_logic;                                        -- chipselect
			SPI_ENET_spi_control_port_address         : out std_logic_vector(2 downto 0);                     -- address
			SPI_ENET_spi_control_port_write           : out std_logic;                                        -- write
			SPI_ENET_spi_control_port_read            : out std_logic;                                        -- read
			SPI_ENET_spi_control_port_readdata        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SPI_ENET_spi_control_port_writedata       : out std_logic_vector(15 downto 0);                    -- writedata
			SPI_ENET_spi_control_port_chipselect      : out std_logic;                                        -- chipselect
			SystemTick_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			SystemTick_s1_write                       : out std_logic;                                        -- write
			SystemTick_s1_readdata                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SystemTick_s1_writedata                   : out std_logic_vector(15 downto 0);                    -- writedata
			SystemTick_s1_chipselect                  : out std_logic                                         -- chipselect
		);
	end component nios_mm_interconnect_0;

	component nios_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                                     : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                         : std_logic_vector(15 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                            : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_write                                           : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                       : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                  : std_logic_vector(17 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                     : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest               : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_ram_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	signal mm_interconnect_0_ram_s1_readdata                               : std_logic_vector(31 downto 0); -- RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	signal mm_interconnect_0_ram_s1_address                                : std_logic_vector(10 downto 0); -- mm_interconnect_0:RAM_s1_address -> RAM:address
	signal mm_interconnect_0_ram_s1_byteenable                             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	signal mm_interconnect_0_ram_s1_write                                  : std_logic;                     -- mm_interconnect_0:RAM_s1_write -> RAM:write
	signal mm_interconnect_0_ram_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	signal mm_interconnect_0_ram_s1_clken                                  : std_logic;                     -- mm_interconnect_0:RAM_s1_clken -> RAM:clken
	signal mm_interconnect_0_gpio_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:GPIO_s1_chipselect -> GPIO:chipselect
	signal mm_interconnect_0_gpio_s1_readdata                              : std_logic_vector(31 downto 0); -- GPIO:readdata -> mm_interconnect_0:GPIO_s1_readdata
	signal mm_interconnect_0_gpio_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:GPIO_s1_address -> GPIO:address
	signal mm_interconnect_0_gpio_s1_write                                 : std_logic;                     -- mm_interconnect_0:GPIO_s1_write -> mm_interconnect_0_gpio_s1_write:in
	signal mm_interconnect_0_gpio_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:GPIO_s1_writedata -> GPIO:writedata
	signal mm_interconnect_0_systemtick_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:SystemTick_s1_chipselect -> SystemTick:chipselect
	signal mm_interconnect_0_systemtick_s1_readdata                        : std_logic_vector(15 downto 0); -- SystemTick:readdata -> mm_interconnect_0:SystemTick_s1_readdata
	signal mm_interconnect_0_systemtick_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SystemTick_s1_address -> SystemTick:address
	signal mm_interconnect_0_systemtick_s1_write                           : std_logic;                     -- mm_interconnect_0:SystemTick_s1_write -> mm_interconnect_0_systemtick_s1_write:in
	signal mm_interconnect_0_systemtick_s1_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:SystemTick_s1_writedata -> SystemTick:writedata
	signal mm_interconnect_0_spi_enet_spi_control_port_chipselect          : std_logic;                     -- mm_interconnect_0:SPI_ENET_spi_control_port_chipselect -> SPI_ENET:spi_select
	signal mm_interconnect_0_spi_enet_spi_control_port_readdata            : std_logic_vector(15 downto 0); -- SPI_ENET:data_to_cpu -> mm_interconnect_0:SPI_ENET_spi_control_port_readdata
	signal mm_interconnect_0_spi_enet_spi_control_port_address             : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SPI_ENET_spi_control_port_address -> SPI_ENET:mem_addr
	signal mm_interconnect_0_spi_enet_spi_control_port_read                : std_logic;                     -- mm_interconnect_0:SPI_ENET_spi_control_port_read -> mm_interconnect_0_spi_enet_spi_control_port_read:in
	signal mm_interconnect_0_spi_enet_spi_control_port_write               : std_logic;                     -- mm_interconnect_0:SPI_ENET_spi_control_port_write -> mm_interconnect_0_spi_enet_spi_control_port_write:in
	signal mm_interconnect_0_spi_enet_spi_control_port_writedata           : std_logic_vector(15 downto 0); -- mm_interconnect_0:SPI_ENET_spi_control_port_writedata -> SPI_ENET:data_from_cpu
	signal mm_interconnect_0_spi_eeprom_spi_control_port_chipselect        : std_logic;                     -- mm_interconnect_0:SPI_EEPROM_spi_control_port_chipselect -> SPI_EEPROM:spi_select
	signal mm_interconnect_0_spi_eeprom_spi_control_port_readdata          : std_logic_vector(15 downto 0); -- SPI_EEPROM:data_to_cpu -> mm_interconnect_0:SPI_EEPROM_spi_control_port_readdata
	signal mm_interconnect_0_spi_eeprom_spi_control_port_address           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SPI_EEPROM_spi_control_port_address -> SPI_EEPROM:mem_addr
	signal mm_interconnect_0_spi_eeprom_spi_control_port_read              : std_logic;                     -- mm_interconnect_0:SPI_EEPROM_spi_control_port_read -> mm_interconnect_0_spi_eeprom_spi_control_port_read:in
	signal mm_interconnect_0_spi_eeprom_spi_control_port_write             : std_logic;                     -- mm_interconnect_0:SPI_EEPROM_spi_control_port_write -> mm_interconnect_0_spi_eeprom_spi_control_port_write:in
	signal mm_interconnect_0_spi_eeprom_spi_control_port_writedata         : std_logic_vector(15 downto 0); -- mm_interconnect_0:SPI_EEPROM_spi_control_port_writedata -> SPI_EEPROM:data_from_cpu
	signal mm_interconnect_0_rom_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:ROM_s1_chipselect -> ROM:chipselect
	signal mm_interconnect_0_rom_s1_readdata                               : std_logic_vector(31 downto 0); -- ROM:readdata -> mm_interconnect_0:ROM_s1_readdata
	signal mm_interconnect_0_rom_s1_debugaccess                            : std_logic;                     -- mm_interconnect_0:ROM_s1_debugaccess -> ROM:debugaccess
	signal mm_interconnect_0_rom_s1_address                                : std_logic_vector(12 downto 0); -- mm_interconnect_0:ROM_s1_address -> ROM:address
	signal mm_interconnect_0_rom_s1_byteenable                             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ROM_s1_byteenable -> ROM:byteenable
	signal mm_interconnect_0_rom_s1_write                                  : std_logic;                     -- mm_interconnect_0:ROM_s1_write -> ROM:write
	signal mm_interconnect_0_rom_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:ROM_s1_writedata -> ROM:writedata
	signal mm_interconnect_0_rom_s1_clken                                  : std_logic;                     -- mm_interconnect_0:ROM_s1_clken -> ROM:clken
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- SPI_ENET:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- SPI_EEPROM:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- SystemTick:irq -> irq_mapper:receiver3_irq
	signal cpu_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [RAM:reset, ROM:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, ROM:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_gpio_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_gpio_s1_write:inv -> GPIO:write_n
	signal mm_interconnect_0_systemtick_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_systemtick_s1_write:inv -> SystemTick:write_n
	signal mm_interconnect_0_spi_enet_spi_control_port_read_ports_inv      : std_logic;                     -- mm_interconnect_0_spi_enet_spi_control_port_read:inv -> SPI_ENET:read_n
	signal mm_interconnect_0_spi_enet_spi_control_port_write_ports_inv     : std_logic;                     -- mm_interconnect_0_spi_enet_spi_control_port_write:inv -> SPI_ENET:write_n
	signal mm_interconnect_0_spi_eeprom_spi_control_port_read_ports_inv    : std_logic;                     -- mm_interconnect_0_spi_eeprom_spi_control_port_read:inv -> SPI_EEPROM:read_n
	signal mm_interconnect_0_spi_eeprom_spi_control_port_write_ports_inv   : std_logic;                     -- mm_interconnect_0_spi_eeprom_spi_control_port_write:inv -> SPI_EEPROM:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, GPIO:reset_n, SPI_EEPROM:reset_n, SPI_ENET:reset_n, SystemTick:reset_n, jtag_uart_0:rst_n]

begin

	cpu : component nios_CPU
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                              --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	gpio : component nios_GPIO
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_gpio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_gpio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_gpio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_gpio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_gpio_s1_readdata,        --                    .readdata
			out_port   => gpio_export                                -- external_connection.export
		);

	ram : component nios_RAM
		port map (
			clk        => clk_clk,                             --   clk1.clk
			address    => mm_interconnect_0_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,  --       .reset_req
			freeze     => '0'                                  -- (terminated)
		);

	rom : component nios_ROM
		port map (
			clk         => clk_clk,                              --   clk1.clk
			address     => mm_interconnect_0_rom_s1_address,     --     s1.address
			debugaccess => mm_interconnect_0_rom_s1_debugaccess, --       .debugaccess
			clken       => mm_interconnect_0_rom_s1_clken,       --       .clken
			chipselect  => mm_interconnect_0_rom_s1_chipselect,  --       .chipselect
			write       => mm_interconnect_0_rom_s1_write,       --       .write
			readdata    => mm_interconnect_0_rom_s1_readdata,    --       .readdata
			writedata   => mm_interconnect_0_rom_s1_writedata,   --       .writedata
			byteenable  => mm_interconnect_0_rom_s1_byteenable,  --       .byteenable
			reset       => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze      => '0'                                   -- (terminated)
		);

	spi_eeprom : component nios_SPI_EEPROM
		port map (
			clk           => clk_clk,                                                       --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                      --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_eeprom_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_eeprom_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_eeprom_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_eeprom_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_eeprom_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_eeprom_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver2_irq,                                      --              irq.irq
			MISO          => spi_eeprom_external_MISO,                                      --         external.export
			MOSI          => spi_eeprom_external_MOSI,                                      --                 .export
			SCLK          => spi_eeprom_external_SCLK,                                      --                 .export
			SS_n          => spi_eeprom_external_SS_n                                       --                 .export
		);

	spi_enet : component nios_SPI_ENET
		port map (
			clk           => clk_clk,                                                     --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                    --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_enet_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_enet_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_enet_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_enet_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_enet_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_enet_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver1_irq,                                    --              irq.irq
			MISO          => spi_enet_external_MISO,                                      --         external.export
			MOSI          => spi_enet_external_MOSI,                                      --                 .export
			SCLK          => spi_enet_external_SCLK,                                      --                 .export
			SS_n          => spi_enet_external_SS_n                                       --                 .export
		);

	systemtick : component nios_SystemTick
		port map (
			clk        => clk_clk,                                         --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			address    => mm_interconnect_0_systemtick_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_systemtick_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_systemtick_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_systemtick_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_systemtick_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                         --   irq.irq
		);

	jtag_uart_0 : component nios_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	mm_interconnect_0 : component nios_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                                     --                       clk_0_clk.clk
			CPU_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                              -- CPU_reset_reset_bridge_in_reset.reset
			CPU_data_master_address                   => cpu_data_master_address,                                     --                 CPU_data_master.address
			CPU_data_master_waitrequest               => cpu_data_master_waitrequest,                                 --                                .waitrequest
			CPU_data_master_byteenable                => cpu_data_master_byteenable,                                  --                                .byteenable
			CPU_data_master_read                      => cpu_data_master_read,                                        --                                .read
			CPU_data_master_readdata                  => cpu_data_master_readdata,                                    --                                .readdata
			CPU_data_master_write                     => cpu_data_master_write,                                       --                                .write
			CPU_data_master_writedata                 => cpu_data_master_writedata,                                   --                                .writedata
			CPU_data_master_debugaccess               => cpu_data_master_debugaccess,                                 --                                .debugaccess
			CPU_instruction_master_address            => cpu_instruction_master_address,                              --          CPU_instruction_master.address
			CPU_instruction_master_waitrequest        => cpu_instruction_master_waitrequest,                          --                                .waitrequest
			CPU_instruction_master_read               => cpu_instruction_master_read,                                 --                                .read
			CPU_instruction_master_readdata           => cpu_instruction_master_readdata,                             --                                .readdata
			CPU_debug_mem_slave_address               => mm_interconnect_0_cpu_debug_mem_slave_address,               --             CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write                 => mm_interconnect_0_cpu_debug_mem_slave_write,                 --                                .write
			CPU_debug_mem_slave_read                  => mm_interconnect_0_cpu_debug_mem_slave_read,                  --                                .read
			CPU_debug_mem_slave_readdata              => mm_interconnect_0_cpu_debug_mem_slave_readdata,              --                                .readdata
			CPU_debug_mem_slave_writedata             => mm_interconnect_0_cpu_debug_mem_slave_writedata,             --                                .writedata
			CPU_debug_mem_slave_byteenable            => mm_interconnect_0_cpu_debug_mem_slave_byteenable,            --                                .byteenable
			CPU_debug_mem_slave_waitrequest           => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,           --                                .waitrequest
			CPU_debug_mem_slave_debugaccess           => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,           --                                .debugaccess
			GPIO_s1_address                           => mm_interconnect_0_gpio_s1_address,                           --                         GPIO_s1.address
			GPIO_s1_write                             => mm_interconnect_0_gpio_s1_write,                             --                                .write
			GPIO_s1_readdata                          => mm_interconnect_0_gpio_s1_readdata,                          --                                .readdata
			GPIO_s1_writedata                         => mm_interconnect_0_gpio_s1_writedata,                         --                                .writedata
			GPIO_s1_chipselect                        => mm_interconnect_0_gpio_s1_chipselect,                        --                                .chipselect
			jtag_uart_0_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --   jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                .write
			jtag_uart_0_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                .read
			jtag_uart_0_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                .readdata
			jtag_uart_0_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                .chipselect
			RAM_s1_address                            => mm_interconnect_0_ram_s1_address,                            --                          RAM_s1.address
			RAM_s1_write                              => mm_interconnect_0_ram_s1_write,                              --                                .write
			RAM_s1_readdata                           => mm_interconnect_0_ram_s1_readdata,                           --                                .readdata
			RAM_s1_writedata                          => mm_interconnect_0_ram_s1_writedata,                          --                                .writedata
			RAM_s1_byteenable                         => mm_interconnect_0_ram_s1_byteenable,                         --                                .byteenable
			RAM_s1_chipselect                         => mm_interconnect_0_ram_s1_chipselect,                         --                                .chipselect
			RAM_s1_clken                              => mm_interconnect_0_ram_s1_clken,                              --                                .clken
			ROM_s1_address                            => mm_interconnect_0_rom_s1_address,                            --                          ROM_s1.address
			ROM_s1_write                              => mm_interconnect_0_rom_s1_write,                              --                                .write
			ROM_s1_readdata                           => mm_interconnect_0_rom_s1_readdata,                           --                                .readdata
			ROM_s1_writedata                          => mm_interconnect_0_rom_s1_writedata,                          --                                .writedata
			ROM_s1_byteenable                         => mm_interconnect_0_rom_s1_byteenable,                         --                                .byteenable
			ROM_s1_chipselect                         => mm_interconnect_0_rom_s1_chipselect,                         --                                .chipselect
			ROM_s1_clken                              => mm_interconnect_0_rom_s1_clken,                              --                                .clken
			ROM_s1_debugaccess                        => mm_interconnect_0_rom_s1_debugaccess,                        --                                .debugaccess
			SPI_EEPROM_spi_control_port_address       => mm_interconnect_0_spi_eeprom_spi_control_port_address,       --     SPI_EEPROM_spi_control_port.address
			SPI_EEPROM_spi_control_port_write         => mm_interconnect_0_spi_eeprom_spi_control_port_write,         --                                .write
			SPI_EEPROM_spi_control_port_read          => mm_interconnect_0_spi_eeprom_spi_control_port_read,          --                                .read
			SPI_EEPROM_spi_control_port_readdata      => mm_interconnect_0_spi_eeprom_spi_control_port_readdata,      --                                .readdata
			SPI_EEPROM_spi_control_port_writedata     => mm_interconnect_0_spi_eeprom_spi_control_port_writedata,     --                                .writedata
			SPI_EEPROM_spi_control_port_chipselect    => mm_interconnect_0_spi_eeprom_spi_control_port_chipselect,    --                                .chipselect
			SPI_ENET_spi_control_port_address         => mm_interconnect_0_spi_enet_spi_control_port_address,         --       SPI_ENET_spi_control_port.address
			SPI_ENET_spi_control_port_write           => mm_interconnect_0_spi_enet_spi_control_port_write,           --                                .write
			SPI_ENET_spi_control_port_read            => mm_interconnect_0_spi_enet_spi_control_port_read,            --                                .read
			SPI_ENET_spi_control_port_readdata        => mm_interconnect_0_spi_enet_spi_control_port_readdata,        --                                .readdata
			SPI_ENET_spi_control_port_writedata       => mm_interconnect_0_spi_enet_spi_control_port_writedata,       --                                .writedata
			SPI_ENET_spi_control_port_chipselect      => mm_interconnect_0_spi_enet_spi_control_port_chipselect,      --                                .chipselect
			SystemTick_s1_address                     => mm_interconnect_0_systemtick_s1_address,                     --                   SystemTick_s1.address
			SystemTick_s1_write                       => mm_interconnect_0_systemtick_s1_write,                       --                                .write
			SystemTick_s1_readdata                    => mm_interconnect_0_systemtick_s1_readdata,                    --                                .readdata
			SystemTick_s1_writedata                   => mm_interconnect_0_systemtick_s1_writedata,                   --                                .writedata
			SystemTick_s1_chipselect                  => mm_interconnect_0_systemtick_s1_chipselect                   --                                .chipselect
		);

	irq_mapper : component nios_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_gpio_s1_write_ports_inv <= not mm_interconnect_0_gpio_s1_write;

	mm_interconnect_0_systemtick_s1_write_ports_inv <= not mm_interconnect_0_systemtick_s1_write;

	mm_interconnect_0_spi_enet_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_enet_spi_control_port_read;

	mm_interconnect_0_spi_enet_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_enet_spi_control_port_write;

	mm_interconnect_0_spi_eeprom_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_eeprom_spi_control_port_read;

	mm_interconnect_0_spi_eeprom_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_eeprom_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios
